$date
	Sat Aug 27 23:49:40 2022
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module fa_tb $end
$var wire 1 ! s $end
$var wire 1 " c $end
$var reg 1 # a $end
$var reg 1 $ b $end
$var reg 1 % cin $end
$scope module fa1 $end
$var wire 1 # a $end
$var wire 1 $ b $end
$var wire 1 % cin $end
$var reg 1 " c $end
$var reg 1 ! s $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0%
0$
0#
0"
0!
$end
#20
1!
1%
#30
1$
0%
#40
1"
0!
1%
#50
0"
1!
1#
0$
0%
#60
1"
0!
1%
#70
1$
0%
#80
1!
1%
